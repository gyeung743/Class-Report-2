module disp_hex_mux (
    input  logic clk, reset,
    input  logic [3:0] hex3, hex2, hex1, hex0, // hex digits
    input  logic [3:0] dp_in,                  // 4 decimal points
    output logic [3:0] an,                     // enable
    output logic [7:0] sseg                    // led segments
);

    // constant declaration
    // refreshing rate around 800 Hz (50 MHz / 2^16)
    localparam N = 18;
    // internal signal declaration
    logic [N-1:0] q_reg;
    logic [N-1:0] q_next;
    logic [3:0] hex_in;
    logic dp;

    // N-bit counter
    always_ff @(posedge clk, posedge reset)
        if (reset)
            q_reg <= 0;
        else
            q_reg <= q_next;

    // next-state logic
    assign q_next = q_reg + 1;

    // 2 MSBs of counter to control 4-to-1 multiplexing and to generate active-low enable signal
    always_comb
        case (q_reg[N-1:N-2])
            2'b00: begin
                an     = 4'b1110;
                hex_in = hex0;
                dp     = dp_in[0];
            end
            2'b01: begin
                an     = 4'b1101;
                hex_in = hex1;
                dp     = dp_in[1];
            end
            2'b10: begin
                an     = 4'b1011;
                hex_in = hex2;
                dp     = dp_in[2];
            end
            default: begin
                an     = 4'b0111;
                hex_in = hex3;
                dp     = dp_in[3];
            end
        endcase

    // hex to seven-segment led display
    always_comb
        case (hex_in)
            4'h0:     sseg[6:0] = 7'b1000000;
            4'h1:     sseg[6:0] = 7'b1111001;
            4'h2:     sseg[6:0] = 7'b0100100;
            4'h3:     sseg[6:0] = 7'b0110000;
            4'h4:     sseg[6:0] = 7'b0011001;
            4'h5:     sseg[6:0] = 7'b0010010;
            4'h6:     sseg[6:0] = 7'b0000010;
            4'h7:     sseg[6:0] = 7'b1111000;
            4'h8:     sseg[6:0] = 7'b0000000;
            4'h9:     sseg[6:0] = 7'b0010000;
            4'hA:     sseg[6:0] = 7'b0001000;
            4'hB:     sseg[6:0] = 7'b0000011;
            4'hC:     sseg[6:0] = 7'b1000110;
            4'hD:     sseg[6:0] = 7'b0100001;
            4'hE:     sseg[6:0] = 7'b0000110;
            default:  sseg[6:0] = 7'b0001110; // 4'hF
        endcase

    assign sseg[7] = dp;

endmodule
